module RegisterFile
(
	input  wire   Clk,
	input  wire   iWE,
	input  wire   [4:0] iWA, iRA1, iRA2,
    input  wire   [31:0] iWD,
    output logic  [31:0] oRD1, oRD2
);

endmodule

