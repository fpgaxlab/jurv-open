module Controller(
   input  wire  [6:0] iOpcode,
   input  wire  [2:0] iFunct3,
   output logic oRegWrite,   
   output riscv_defs::t_imm oImmType
);

endmodule

